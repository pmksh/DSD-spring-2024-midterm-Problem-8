library verilog;
use verilog.vl_types.all;
entity Parking_test_4 is
end Parking_test_4;
