library verilog;
use verilog.vl_types.all;
entity Parking_test_2 is
end Parking_test_2;
