library verilog;
use verilog.vl_types.all;
entity Parking_test is
end Parking_test;
