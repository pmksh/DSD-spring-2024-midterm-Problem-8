library verilog;
use verilog.vl_types.all;
entity Parking_test_3 is
end Parking_test_3;
